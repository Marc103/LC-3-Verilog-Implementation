module BUS_DRIVER(input [15:0] MARMUX_OUT,
                  input [15:0] PC_OUT,
                  input [15:0]
                   output [15:0] BUS);
    reg [15:0] Result;       

...